library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity AIRFRYER is
end AIRFRYER;

architecture Behavioral of AIRFRYER is
   signal boton_sync: std_logic;
   signal boton_edge: std_logic;
begin


end Behavioral;
